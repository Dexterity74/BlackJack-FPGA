/*	file name: card.svh
	Authors: Justin Negron and Richard Osborn
	created: 08/06/21
	team name: POWER_OF_TWO

	signal that represents card values
*/

//custom signal type
typedef logic [3:0] card;
