/*	file name: dealerAI
	Authors: Justin Negron and Richard Osborn
	created: 07/30/21
	team name: POWER_OF_TWO

	describes a hand of cards
	represents the sum of all the cards in the player's hand.
	must cover [0, 30] //worst hand is three 10s.
	2 ^ 5 = 32

*/

typedef logic [4 : 0] hand;
