/*	file name: dealerAI
	Authors: Justin Negron and Richard Osborn
	created: 07/30/21
	team name: POWER_OF_TWO
*/

//custom signal type
//package blackjack;
typedef enum logic [2:0] {NONE, HIT, STAND, DOUBLE} gameCommand;
//endpackage