/*	file name: card.svh
	Authors: Justin Negron and Richard Osborn
	created: 08/06/21
	team name: POWER_OF_TWO

	signal that represents card values
*/

//custom signal type
`define card logic [3:0]
`define MAX_CARDS 5
`define CARD_WIDTH 4
//typedef logic [3:0] card;
