/*	file name: card.svh
	Authors: Justin Negron and Richard Osborn
	created: 08/06/21
	team name: POWER_OF_TWO

	signal that represents card values
*/

//custom signal type
`define card logic [3:0]
`define HAND_OF_5_CARDS logic [3:0] [4:0] //5 cards of 4 bits
`define MAX_CARDS 5
//typedef logic [3:0] card;
