/*	file name: blackjackGame
	Authors: Justin Negron and Richard Osborn
	created: 07/30/21
	team name: POWER_OF_TWO
*/

module blackjackGame
	(
		input  logic 	      clk,
		input  logic 	      reset,
		input  logic 		  hit, stand,
	);
endmodule