/*	file name: dealerAI
	Authors: Justin Negron and Richard Osborn
	created: 07/30/21
	team name: POWER_OF_TWO

	describes a hand of cards

*/

//wtf??? why doesn't this work?


package blackjack;

typedef logic [4 : 0] hand;
endpackage